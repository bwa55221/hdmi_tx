LIBRARY ieee;
USE ieee.std_logic_1164.all;

package custom_pkg is
    type iic_data_array is array(0 to 1) of std_logic_vector(7 downto 0);
end custom_pkg;

package body custom_pkg is

end custom_pkg;